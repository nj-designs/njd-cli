//------------------------------------------------------------------
//-- Hello world example
//-- Turn on all the leds
//-- This example has been tested on the following boards:
//--   * Lattice icestick
//--   * Icezum alhambra (https://github.com/FPGAwars/icezum)
//------------------------------------------------------------------

module led_adder(output wire LED0,
                 output wire LED1);

assign LED0 = 1'b1;
assign LED1 = 1'b1;

endmodule
